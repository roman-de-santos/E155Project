`timescale 1ns / 1ps

module Data_Slow_to_Fast_tb;

    // =========================================================================
    // 1. Parameters & Signals
    // =========================================================================
    parameter WIDTH = 16;
    
    // Simulation Clocks
    logic Clk_Fast = 0; // 6 MHz (DSP System Clock)
    logic Clk_Slow = 0; // ~1.41 MHz (I2S Bit Clock)
    
    // Control Signals
    logic Rst = 1;
    
    // Slow Domain Inputs (Drivers)
    logic [WIDTH-1:0] Data_In_Slow;
    logic             Valid_In_Slow;
    
    // Fast Domain Outputs (Monitors)
    logic [WIDTH-1:0] Data_Out_Fast;
    logic             Valid_Out_Fast;

    // Test Variables
    logic [WIDTH-1:0] expected_data;
    integer error_count = 0;
    integer transaction_count = 0;

    // =========================================================================
    // 2. DUT Instantiation
    // =========================================================================
    Data_Slow_to_Fast #(
        .WIDTH(WIDTH)
    ) DUT (
        .Clk_Fast(Clk_Fast),
        .Rst(Rst),
        .Data_In_Slow(Data_In_Slow),
        .Valid_In_Slow(Valid_In_Slow),
        .Data_Out_Fast(Data_Out_Fast),
        .Valid_Out_Fast(Valid_Out_Fast)
    );

    // =========================================================================
    // 3. Clock Generation
    // =========================================================================
    
    // 6 MHz Fast Clock -> Period approx 166.6 ns
    // Half period = 83.3 ns
    always #83.3 Clk_Fast = ~Clk_Fast; 

    // 1.41 MHz Slow Clock -> Period approx 709 ns
    // Half period = 354.5 ns
    // We add a tiny offset to make it asynchronous (real world simulation)
    always #354.5 Clk_Slow = ~Clk_Slow; 

    // =========================================================================
    // 4. Test Sequence
    // =========================================================================
    initial begin
        $display("=== Starting Slow to Fast CDC Testbench ===");
        $display("Ref: Fast Clock = 6MHz, Slow Clock = 1.41MHz");
        
        // Initialize
        Rst = 1;
        Valid_In_Slow = 0;
        Data_In_Slow = 0;
        
        // Apply Reset
        #500;
        @(posedge Clk_Fast);
        Rst = 0; // Active High Reset in your module? (Check your module, I assumed active high)
                 // NOTE: Your top.sv uses ~rst (Active Low button), but typically internal resets are active high or low.
                 // In the module code provided earlier: "if (Rst)..." implies Active High.
        
        $display("Reset Released");
        #200;

        // --- Transaction Loop ---
        repeat (10) begin
            // 1. Generate Random Data
            expected_data = $urandom();
            
            // 2. Drive Data in SLOW Domain
            // We align to the Slow Clock to mimic I2S Rx behavior
            @(posedge Clk_Slow);
            Data_In_Slow  <= expected_data;
            Valid_In_Slow <= 1'b1; 
            
            // Hold the signal HIGH for one full slow cycle (mimicking the WS edge logic)
            // Note: In reality, WS might be high for 16 slow clocks, but a 1-cycle pulse
            // generated by edge detection logic in top.sv is what enters here.
            @(posedge Clk_Slow); 
            Valid_In_Slow <= 1'b0;
            
            // 3. Monitor FAST Domain Output
            // The Fast clock runs 4x faster. It should catch this.
            
            fork
                begin
                    // Wait for the pulse in Fast Domain
                    @(posedge Valid_Out_Fast); 
                end
                begin
                    // Timeout watchdog (approx 5 slow cycles)
                    #3500; 
                    $display("ERROR: Timeout waiting for data transfer!");
                    $stop;
                end
            join_any
            disable fork;

            // 4. Check Data
            // We check slightly after the edge to ensure stability
            #1; 
            if (Data_Out_Fast === expected_data) begin
                $display("[PASS] Time: %0t | Sent: 0x%h | Received: 0x%h", $time, expected_data, Data_Out_Fast);
            end else begin
                $display("[FAIL] Time: %0t | Sent: 0x%h | Received: 0x%h", $time, expected_data, Data_Out_Fast);
                error_count++;
            end

            // 5. Check for "Double Trigger" (Crucial for Slow->Fast)
            // Ensure Valid_Out_Fast goes LOW immediately after 1 cycle.
            @(posedge Clk_Fast);
            if (Valid_Out_Fast == 1'b1) begin
                $display("[FAIL] Valid_Out_Fast stuck HIGH for more than 1 cycle!");
                error_count++;
            end

            transaction_count++;
            
            // Random Delay before next packet
            repeat ($urandom_range(2, 5)) @(posedge Clk_Slow);
        end

        // --- Final Report ---
        #1000;
        if (error_count == 0)
            $display("=== TEST PASSED: %0d Transactions Successful ===", transaction_count);
        else
            $display("=== TEST FAILED: %0d Errors Detected ===", error_count);
        
        $finish;
    end

endmodule